`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/27/2019 12:27:05 PM
// Design Name: 
// Module Name: q6tic
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module q6tic(v11,v12,v13,v21,v22,v23,v31,v32,v33,p,win);
input [2:0]v11,v12,v13,v21,v22,v23,v31,v32,v33;//data for 9 tic tac toe blocks
output win;//1 indicates player can win
reg win;
input p;//indicates which player's turn
always@(*)
begin
if (p==1)
begin
if((v11==3 && v12==3 && (v13!=0 && v13!=3)) ||
(v11==3 && v13==3 && (v12!=0 && v12!=3))||
(v13==3 && v12==3 && (v11!=0 && v11!=3))||
(v21==3 && v22==3 && (v23!=0 && v23!=3))||
(v23==3 && v22==3 && (v21!=0 && v21!=3))||
(v23==3 && v21==3 && (v22!=0 && v22!=3))||
(v31==3 && v32==3 && (v33!=0 && v33!=3))||
(v33==3 && v32==3 && (v31!=0 && v31!=3))||
(v11==3 && v21==3 && (v31!=0 && v31!=3))||
(v11==3 && v31==3 && (v21!=0 && v21!=3))||
(v21==3 && v31==3 && (v11!=0 && v11!=3))||
(v12==3 && v22==3 && (v32!=0 && v32!=3))||
(v22==3 && v23==3 && (v12!=0 && v12!=3))||
(v32==3 && v21==3 && (v22!=0 && v22!=3))||
(v13==3 && v23==3 && (v33!=0 && v33!=3))||
(v23==3 && v33==3 && (v13!=0 && v13!=3))||
(v33==3 && v13==3 && (v22!=0 && v22!=3))||
(v11==3 && v22==3 && (v33!=0 && v33!=3))||
(v33==3 && v11==3 && (v22!=0 && v22!=3))||
(v22==3 && v33==3 && (v11!=0 && v11!=3))||
(v13==3 && v31==3 && (v22!=0 && v22!=3))||
(v22==3 && v13==3 && (v31!=0 && v31!=3))||
(v31==3 && v22==3 && (v13!=0 && v13!=3)))//checking for all cases for player 1
win=1;
end
if(p==0)
begin
if((v11==3 && v12==3 && (v13!=0 && v13!=3)) ||
(v11==0 && v13==0 && (v12!=0 && v12!=3))||
(v13==0 && v12==0 && (v11!=0 && v11!=3))||
(v21==0 && v22==0 && (v23!=0 && v23!=3))||
(v23==0 && v22==0 && (v21!=0 && v21!=3))||
(v23==0 && v21==0 && (v22!=0 && v22!=3))||
(v31==0 && v32==0 && (v33!=0 && v33!=3))||
(v33==0 && v32==0 && (v31!=0 && v31!=3))||
(v11==0 && v21==0 && (v31!=0 && v31!=3))||
(v11==0 && v31==0 && (v21!=0 && v21!=3))||
(v21==0 && v31==0 && (v11!=0 && v11!=3))||
(v12==0 && v22==0 && (v32!=0 && v32!=3))||
(v22==0 && v23==0 && (v12!=0 && v12!=3))||
(v32==0 && v21==0 && (v22!=0 && v22!=3))||
(v13==0 && v23==0 && (v33!=0 && v33!=3))||
(v23==0 && v33==0 && (v13!=0 && v13!=3))||
(v33==0 && v13==0 && (v22!=0 && v22!=3))||
(v33==0 && v13==0 && (v22!=0 && v22!=3))||
(v11==0 && v22==0 && (v33!=0 && v33!=3))||
(v33==0 && v11==0 && (v22!=0 && v22!=3))||
(v22==0 && v33==0 && (v11!=0 && v11!=3))||
(v13==0 && v31==0 && (v22!=0 && v22!=3))||
(v22==0 && v13==0 && (v31!=0 && v31!=3))||
(v31==0 && v22==0 && (v13!=0 && v13!=3)))//checking for all cases for player 2
win=1;
end
if(win!=1)
begin
win=0;
end
end


endmodule

